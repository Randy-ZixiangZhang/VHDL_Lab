----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:16:40 02/02/2022 
-- Design Name: 
-- Module Name:    mux4x1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux4x1 is

	port(S: in STD_LOGIC_VECTOR(1 downto 0);
		  D0 : in  STD_LOGIC_VECTOR (15 downto 0);
		  D1 : in  STD_LOGIC_VECTOR (15 downto 0);
		  D2 : in  STD_LOGIC_VECTOR (15 downto 0);
		  D3 : in  STD_LOGIC_VECTOR (15 downto 0);
		  O: out STD_LOGIC_VECTOR (15 downto 0));


end mux4x1;

architecture Behavioral of mux4x1 is

begin

	process(S,D0,D1,D2,D3) is
	begin
		case S is
			when "00" =>
				O <= D0;
			when "01" =>
				O <= D1;
			when "10" =>
				O <= D2;
			when "11" =>
				O <= D3;
			when others =>
				O <= "XXXXXXXXXXXXXXXX"; --must use "", error using ''
		end case;
	end process;

end Behavioral;

